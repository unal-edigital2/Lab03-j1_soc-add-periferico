module display( input [7:0] bcd, output [6:0] sseg_d1, output [6:0] sseg_d2);

// tambien colocar las señales de control que hacen falta en el bloque ejemplo clk
//colocar aca el codigo que hace falta y que ya lo tienen de los laboratorios anteriores

endmodule
